module Processor ()


endmodule
